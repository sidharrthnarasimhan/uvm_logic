interface halfadder_intf;
    logic sig_clock;
    logic sig_in_a;
    logic sig_in_b;
    logic sig_reset;
    logic sig_carry;
    logic sig_sum;
endinterface: halfadder_intf