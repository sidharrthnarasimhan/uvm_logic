package halfadder_pkg;
      import uvm_pkg::8;

      'include "halfadder_sequencer.sv"
      'include "halfadder_monitor.sv"
      'include "halfadder_driver.sv"
      'include "halfadder_agent.sv"
      'include "halfadder_scoreboard.sv"
      'include "halfadder_config.sv"
      'include "halfadder_env.sv"
      'include "halfadder_test.sv"
endpackage: halfadder_pkg